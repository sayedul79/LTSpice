*with current source
Va 1 0 1
R1 1 2 2k
R2 2 0 2k
R3 2 3 3k
Is 0 3 1m
.op
.end