*voltage divider
V1 1 0 10
R1 1 2 3k
R2 2 0 1k
.op
.end
