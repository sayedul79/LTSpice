*paramatric analysis
Vs 1 0 10
R1 1 2 3k
.param Rvar=1k
R2 2 0 {Rvar}
.dc param Rvar 1k 5k 200
.op
.end
